library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;


entity MemInst is
    Port ( address : in  STD_LOGIC_VECTOR (31 downto 0);
           Instr : out  STD_LOGIC_VECTOR (31 downto 0));
end MemInst;


architecture Behavioral of MemInst is

	type ARRAY_256 is ARRAY (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
	signal MemContent: ARRAY_256 :=	(	
				X"20070040",X"20080048",X"20090060",X"8cea0000",
				X"71072802",X"70C72802",X"71284002",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				x"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000",
				X"00000000",X"00000000",X"00000000",X"00000000");	
	begin

	Instr <= MemContent(to_integer(unsigned(address(31 downto 2))));

end Behavioral;

